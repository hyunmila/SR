//`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////////
//// Company: 
//// Engineer: 
//// 
//// Create Date: 03/07/2023 10:59:12 AM
//// Design Name: 
//// Module Name: linia_opozniajaca
//// Project Name: 
//// Target Devices: 
//// Tool Versions: 
//// Description: 
//// 
//// Dependencies: 
//// 
//// Revision:
//// Revision 0.01 - File Created
//// Additional Comments:
//// 
////////////////////////////////////////////////////////////////////////////////////


//module linia_opozniajaca #
//(
//    parameter N = 1,
//    parameter DELAY = 1
//)
//(
//    input clk,
//    input ce,
//    input idata,
//    output odata
//);
//wire [N-1:0] tdata [DELAY:0];
//genvar i;

//generate
//    if (DELAY == 0)
//    begin
//        assign odata = idata;
//    end
//    if (DELAY > 0)
//    begin
//        for(i=0; i<DELAY; i++)
//        begin
//            DELAY++;
//        end
//    end
//endgenerate

//endmodule


//module one_delay #
//(
//    parameter N = 1
//)
//(
//    input clk,
//    input ce,
//    input d,
//    output [3:0]q
//);
//endmodule